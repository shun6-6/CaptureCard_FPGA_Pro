`define VIVADO